// MU0 ALU design 
// P W Nutter (based on a design by Jeff Pepper)
// Date 7/7/2021

// Do not touch the following line it is required for simulation 
`timescale 1ns/100ps
`default_nettype none

// module header

module MU0_Alu (
               input  wire [15:0]  X, 
               input  wire [15:0]  Y, 
               input  wire [1:0]   M, 
               output reg  [15:0]  Q
	       );

// behavioural description for the ALU







endmodule 

// for simulation purposes, do not delete
`default_nettype wire
